`timescale 1ns/100ps
`include "sar_logic.v"

module tb_sar_logic;

reg rest,clk,comp,ena;
wire []


initial
	begin

	

	end